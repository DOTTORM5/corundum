module packet_transmitter #(
) (
);


memory_fetcher # (

) memory_fetcher_i (

);

packet_builder #(

) packet_builder_i (
    
);


endmodule