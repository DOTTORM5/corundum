module traffic_manager #(
) (
);

filter #(

) filer_i (

);


parser #( 

) parser_i (

);

rule_match_engine #(

) rule_match_engine_i (

);



endmodule