module low_latency_logic #(
) (
);

traffic_manager #(

) traffic_manager_i (

);

packet_transmitter #(

) packet_transmitter_i (

);




endmodule
