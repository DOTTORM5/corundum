`timescale 1ns/1ps


module matcher #(
    parameter AXIS_DATA_WIDTH = 512
) (
    
);
    
endmodule