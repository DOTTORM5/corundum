module packet_builder #(
) (
); 
endmodule